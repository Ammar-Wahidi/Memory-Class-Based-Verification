package Memory_package;

`include "Memory_transaction_class.svh"
`include "Memory_sequencer_class.svh"
`include "Memory_driver_class.svh"
`include "Memory_monitor.svh"
`include "Memory_subscriber_class.svh"
`include "Memory_scoreboard.svh"
`include "Memory_env_class.svh"

endpackage
